package fft_len is
constant LOG2_FFT_LEN : integer := 6;
constant FFT_LEN      : integer := 2 ** LOG2_FFT_LEN;
constant ICPX_WIDTH : integer := 16;
end fft_len;
