package fft_len is
constant LOG2_FFT_LEN : integer := 5;
end fft_len;
