package fft_len is
constant LOG2_FFT_LEN : integer := 9;
end fft_len;
