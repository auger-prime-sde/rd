--- AUGER radio extension FPGA toplevel design

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity top is
  generic (
    -- Number of data bits from the ADC channels
    g_ADC_BITS : natural := 12;
    -- ADC interface width
    g_ADC_DRIVER_BITS : natural := 14;
    -- Number of bits in index counters (11 gives 2048 samples stored)
    g_BUFFER_INDEXSIZE : natural := 11;
    -- Number of bits in serial words
    g_UART_WORDSIZE : natural := 7  );
  port (
    dataIn : in std_logic_vector (g_ADC_DRIVER_BITS-1 downto 0);
    dataOvIn : in std_logic;
    clk : in std_logic;
    rst : in std_logic;
    trigger : in std_logic;
    i_start_transfer : in std_logic;
    o_data : out std_logic);
end top;

architecture behaviour of top is
  constant c_SAMPLE_WIDTH : natural := g_ADC_BITS+1;
  constant c_STORAGE_WIDTH : natural := 2*c_SAMPLE_WIDTH;
  constant c_CLOCK_DIVIDER : natural := 1736;
  constant c_CLOCK_SIZE    : natural := 11;
  constant c_ADC_DRIVER_WIDTH : natural := g_ADC_DRIVER_BITS+1;
  constant c_ADC_DRIVER_OUTPUT_WIDTH : natural := 2*c_ADC_DRIVER_WIDTH;

  signal adc_input_bus : std_logic_vector(c_ADC_DRIVER_WIDTH-1 downto 0);
  signal adc_data : std_logic_vector(c_ADC_DRIVER_OUTPUT_WIDTH-1 downto 0);
  signal adc_data_selected : std_logic_vector(c_STORAGE_WIDTH-1 downto 0);
  signal data_output_bus : std_logic_vector(c_STORAGE_WIDTH-1 downto 0);

  signal buffer_write_en : std_logic;
  signal clk_intern : std_logic;
  signal clk_uart : std_logic;
  signal write_address : std_logic_vector(g_BUFFER_INDEXSIZE-1 downto 0);
  signal read_address : std_logic_vector(g_BUFFER_INDEXSIZE-1 downto 0);
  signal read_set_address : std_logic_vector(g_BUFFER_INDEXSIZE-1 downto 0);

  signal write_trigger_done : std_logic;
  signal write_arm : std_logic;

  signal uart_ready : std_logic;
  signal uart_dataready : std_logic;

  component adc_driver
    port (
      clkin: in  std_logic; reset: in  std_logic; sclk: out  std_logic;
      datain: in  std_logic_vector(c_ADC_DRIVER_WIDTH-1 downto 0);
      q: out  std_logic_vector(c_ADC_DRIVER_OUTPUT_WIDTH-1 downto 0)
    );
  end component;

  component data_buffer
    generic (g_DATA_WIDTH, g_ADDRESS_WIDTH : natural);
    port (
      i_wclk : in std_logic;
      i_we : in std_logic;
      i_waddr : in std_logic_vector(g_BUFFER_INDEXSIZE-1 downto 0);
      i_wdata : in std_logic_vector(c_STORAGE_WIDTH-1 downto 0);
      i_rclk : in std_logic;
      i_re: in std_logic;
      i_raddr : in std_logic_vector(g_BUFFER_INDEXSIZE-1 downto 0);
      o_rdata : out std_logic_vector(c_STORAGE_WIDTH-1 downto 0)
    );
  end component;

  component simple_counter
    generic ( g_SIZE : natural );
    port (
      i_clk: in std_logic;
      o_q: out std_logic_vector(g_BUFFER_INDEXSIZE-1 downto 0)
    );
  end component;

  --component settable_counter
  --  generic ( g_SIZE : natural );
  --  port (
  --    i_en     : in std_logic;
  --    i_clk    : in std_logic;
  --    i_set    : in std_logic;
  --    i_data   : in std_logic_vector(g_BUFFER_INDEXSIZE-1 downto 0);
  --    o_data   : out std_logic_vector(g_BUFFER_INDEXSIZE-1 downto 0)
  --  );
  --end component;

  component uart_expander
    generic (g_WORDSIZE: natural; g_WORDCOUNT : natural);
    port (
      i_data      : in std_logic_vector(g_WORDCOUNT*g_WORDSIZE-1 downto 0);
      i_dataready : in std_logic;
      i_clk       : in std_logic;
      o_data      : out std_logic;
      o_ready     : out std_logic
    );
  end component;

  component write_controller
    generic (g_ADDRESS_BITS : natural; g_START_OFFSET : natural);
    port (
      i_clk          : in std_logic;
      i_trigger      : in std_logic;
      i_curr_addr    : in std_logic_vector(g_ADDRESS_BITS-1 downto 0);
      i_arm          : in std_logic;
      o_write_en     : out std_logic;
      o_trigger_done : out std_logic;
      o_start_addr   : out std_logic_vector(g_ADDRESS_BITS-1 downto 0)
    );
  end component;

  component readout_controller
    generic (g_ADDRESS_BITS : natural);
    port (
      i_clk          : in std_logic;
      i_trigger_done : in std_logic;
      i_start_addr   : in std_logic_vector(g_ADDRESS_BITS-1 downto 0);
      o_arm          : out std_logic := '1';
      o_read_enable  : out std_logic := '1';
      o_read_addr    : out std_logic_vector(g_ADDRESS_BITS-1 downto 0);
      i_word_ready   : in std_logic;
      o_tx_enable    : out std_logic := '0';
      o_tx_ready     : out std_logic := '1';
      i_tx_start     : in std_logic
    );
  end component;

  component clock_divider
    generic (g_SIZE: natural);
    port (
      i_clk     : in std_logic := '0';
      o_clk     : out std_logic := '0';
      i_ratio   : in std_logic_vector(g_SIZE-1 downto 0)
    );
   end component;
begin

  adc_input_bus <= dataOvIn & dataIn;

adc_driver_1 : adc_driver
  port map (
    clkin => clk,
    reset => rst,
    sclk => clk_intern,
    datain =>  adc_input_bus,
    q => adc_data);

  adc_data_selected <=
    adc_data(c_ADC_DRIVER_OUTPUT_WIDTH-1 downto c_ADC_DRIVER_OUTPUT_WIDTH-g_ADC_BITS-1) &
    adc_data(c_ADC_DRIVER_OUTPUT_WIDTH/2-1 downto g_ADC_DRIVER_BITS - g_ADC_BITS);


write_index_counter : simple_counter
  generic map (g_SIZE => g_BUFFER_INDEXSIZE)
  port map (
    i_clk => clk_intern,
    o_q => write_address);

--read_index_counter : settable_counter
--  generic map (g_SIZE => g_BUFFER_INDEXSIZE)
--  port map (
--    i_clk => clk_intern,
--  o_data => read_address,
--  i_en => '1',
--  i_set => '0',
-- i_data => read_set_address);

data_buffer_1 : data_buffer
  generic map (g_ADDRESS_WIDTH => g_BUFFER_INDEXSIZE, g_DATA_WIDTH => c_STORAGE_WIDTH)
  port map (
    i_wclk => clk_intern,
    i_we => buffer_write_en,
    i_waddr => write_address,
    i_rclk => clk_intern,
    i_re => '1',
    i_raddr => read_address,
    i_wdata => adc_data_selected,
    o_rdata => data_output_bus);

uart_1 : uart_expander
  generic map (g_WORDSIZE => g_UART_WORDSIZE, g_WORDCOUNT => 4)
  port map (
    -- TODO: do this more generic:
    i_data(12 downto 0)   => data_output_bus(12 downto 0),
    i_data(26 downto 14)  => data_output_bus(25 downto 13),
    i_data(13)            => '0',
    i_data(27)            => '0',
    i_dataready => uart_dataready,
    i_clk       => clk_uart,
    o_data      => o_data,
    o_ready     => uart_ready
    );



--  o_led <= data_output_bus(0);

write_controller_1 : write_controller
  generic map (g_ADDRESS_BITS => g_BUFFER_INDEXSIZE, g_START_OFFSET => 2047)
  port map (
    i_clk => clk_intern,
    i_trigger => trigger,
    i_curr_addr => write_address,
    i_arm => write_arm,
    o_write_en => buffer_write_en,
    o_start_addr => read_set_address,
    o_trigger_done => open
    );

  readout_controller_1 : readout_controller
    generic map (g_ADDRESS_BITS => g_BUFFER_INDEXSIZE)
    port map (
      i_clk => clk_uart,
      i_trigger_done => write_trigger_done,
      i_start_addr   => read_set_address,
      o_arm          => write_arm,
      o_read_enable  => open,
      o_read_addr    => open,
      i_word_ready   => uart_ready,
      o_tx_enable    => uart_dataready,
      o_tx_ready     => open,
      i_tx_start     => i_start_transfer
   );

  clock_divider_1 : clock_divider
    generic map (g_SIZE => c_CLOCK_SIZE)
    port map (
      i_clk => clk_intern,
      o_clk => clk_uart,
      i_ratio => std_logic_vector(to_unsigned(c_CLOCK_DIVIDER, c_CLOCK_SIZE))
    );

end;
